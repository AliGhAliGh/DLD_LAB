module PWM(clk, rst, inp);
input[7:0] inp;
endmodule